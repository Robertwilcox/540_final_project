/*
 * Authors: Ibrahim Binmahfood, Mohamed Gnedi
 * ECE540, Kravitz
 * Project 2, Character ROM - rtl module
 * 11/18/2023
 *
 * Platform: RVfpga on Boolean Board
 * Description: This module below by default outputs an 8x8 bitmap of 40 ASCII
 * characters. The CLK will be connected via the 25.20 MHz pixel clock. The 8x8
 * bitmaps were originally from: 
 *
 * https://github.com/dhepper/font8x8/blob/master/font8x8_basic.h
 *
 */

module CHAR_ROM #(parameter SIZE = 8, parameter addr_width = 8) (
    input wire logic [addr_width-1:0] address,   // 3-bit address input
	input wire logic CLK,
    output logic [0:SIZE-1] data [0:SIZE-1] // 8-bit data output
);
									
// Declare the ROM content using an initial block
	always_ff @(posedge CLK) begin
		case (address)
//====================================================================================================
// characters || address: [20-23]
//====================================================================================================
			8'h20: data <= {{8'h00}, { 8'h00}, { 8'h00}, { 8'h00}, { 8'h00}, { 8'h00}, { 8'h00}, { 8'h00}}; // space
			8'h21: data <= {{8'h18}, { 8'h3C}, { 8'h3C}, { 8'h18}, { 8'h18}, { 8'h00}, { 8'h18}, { 8'h00}}; // !
			8'h22: data <= {{8'h36}, { 8'h36}, { 8'h00}, { 8'h00}, { 8'h00}, { 8'h00}, { 8'h00}, { 8'h00}}; // "
			8'h23: data <= {{8'h36}, { 8'h36}, { 8'h7F}, { 8'h36}, { 8'h7F}, { 8'h36}, { 8'h36}, { 8'h00}}; // #

//====================================================================================================
// * Numbers {0-9} || address: [30-39]
//====================================================================================================
			8'h30: data <= {{8'h3E}, { 8'h63}, { 8'h73}, { 8'h7B}, { 8'h6F}, { 8'h67}, { 8'h3E}, { 8'h00}}; // 0
			8'h31: data <= {{8'h0C}, { 8'h0E}, { 8'h0C}, { 8'h0C}, { 8'h0C}, { 8'h0C}, { 8'h3F}, { 8'h00}}; // 1
			8'h32: data <= {{8'h1E}, { 8'h33}, { 8'h30}, { 8'h1C}, { 8'h06}, { 8'h33}, { 8'h3F}, { 8'h00}}; // 2
			8'h33: data <= {{8'h1E}, { 8'h33}, { 8'h30}, { 8'h1C}, { 8'h30}, { 8'h33}, { 8'h1E}, { 8'h00}}; // 3
			8'h34: data <= {{8'h38}, { 8'h3C}, { 8'h36}, { 8'h33}, { 8'h7F}, { 8'h30}, { 8'h78}, { 8'h00}}; // 4
			8'h35: data <= {{8'h3F}, { 8'h03}, { 8'h1F}, { 8'h30}, { 8'h30}, { 8'h33}, { 8'h1E}, { 8'h00}}; // 5
			8'h36: data <= {{8'h1C}, { 8'h06}, { 8'h03}, { 8'h1F}, { 8'h33}, { 8'h33}, { 8'h1E}, { 8'h00}}; // 6
			8'h37: data <= {{8'h3F}, { 8'h33}, { 8'h30}, { 8'h18}, { 8'h0C}, { 8'h0C}, { 8'h0C}, { 8'h00}}; // 7
			8'h38: data <= {{8'h1E}, { 8'h33}, { 8'h33}, { 8'h1E}, { 8'h33}, { 8'h33}, { 8'h1E}, { 8'h00}}; // 8
			8'h39: data <= {{8'h1E}, { 8'h33}, { 8'h33}, { 8'h3E}, { 8'h30}, { 8'h18}, { 8'h0E}, { 8'h00}}; // 9
			
//====================================================================================================
// * Letters {a-z} || address: [61-7A]
//====================================================================================================			
			8'h61: data <= {{8'h00}, { 8'h00}, { 8'h1E}, { 8'h30}, { 8'h3E}, { 8'h33}, { 8'h6E}, { 8'h00}}; // a
			8'h62: data <= {{8'h07}, { 8'h06}, { 8'h06}, { 8'h3E}, { 8'h66}, { 8'h66}, { 8'h3B}, { 8'h00}}; // b
			8'h63: data <= {{8'h00}, { 8'h00}, { 8'h1E}, { 8'h33}, { 8'h03}, { 8'h33}, { 8'h1E}, { 8'h00}}; // c
			8'h64: data <= {{8'h38}, { 8'h30}, { 8'h30}, { 8'h3e}, { 8'h33}, { 8'h33}, { 8'h6E}, { 8'h00}}; // d
			8'h65: data <= {{8'h00}, { 8'h00}, { 8'h1E}, { 8'h33}, { 8'h3f}, { 8'h03}, { 8'h1E}, { 8'h00}}; // e
			8'h66: data <= {{8'h1C}, { 8'h36}, { 8'h06}, { 8'h0f}, { 8'h06}, { 8'h06}, { 8'h0F}, { 8'h00}}; // f
			8'h67: data <= {{8'h00}, { 8'h00}, { 8'h6E}, { 8'h33}, { 8'h33}, { 8'h3E}, { 8'h30}, { 8'h1F}}; // g
			8'h68: data <= {{8'h07}, { 8'h06}, { 8'h36}, { 8'h6E}, { 8'h66}, { 8'h66}, { 8'h67}, { 8'h00}}; // h
			8'h69: data <= {{8'h0C}, { 8'h00}, { 8'h0E}, { 8'h0C}, { 8'h0C}, { 8'h0C}, { 8'h1E}, { 8'h00}}; // i
			8'h6A: data <= {{8'h30}, { 8'h00}, { 8'h30}, { 8'h30}, { 8'h30}, { 8'h33}, { 8'h33}, { 8'h1E}}; // j
			8'h6B: data <= {{8'h07}, { 8'h06}, { 8'h66}, { 8'h36}, { 8'h1E}, { 8'h36}, { 8'h67}, { 8'h00}}; // k
			8'h6C: data <= {{8'h0E}, { 8'h0C}, { 8'h0C}, { 8'h0C}, { 8'h0C}, { 8'h0C}, { 8'h1E}, { 8'h00}}; // l
			8'h6D: data <= {{8'h00}, { 8'h00}, { 8'h33}, { 8'h7F}, { 8'h7F}, { 8'h6B}, { 8'h63}, { 8'h00}}; // m
			8'h6E: data <= {{8'h00}, { 8'h00}, { 8'h1F}, { 8'h33}, { 8'h33}, { 8'h33}, { 8'h33}, { 8'h00}}; // n
			8'h6F: data <= {{8'h00}, { 8'h00}, { 8'h1E}, { 8'h33}, { 8'h33}, { 8'h33}, { 8'h1E}, { 8'h00}}; // o
			8'h70: data <= {{8'h00}, { 8'h00}, { 8'h3B}, { 8'h66}, { 8'h66}, { 8'h3E}, { 8'h06}, { 8'h0F}}; // p
			8'h71: data <= {{8'h00}, { 8'h00}, { 8'h6E}, { 8'h33}, { 8'h33}, { 8'h3E}, { 8'h30}, { 8'h78}}; // q
			8'h72: data <= {{8'h00}, { 8'h00}, { 8'h3B}, { 8'h6E}, { 8'h66}, { 8'h06}, { 8'h0F}, { 8'h00}}; // r
			8'h73: data <= {{8'h00}, { 8'h00}, { 8'h3E}, { 8'h03}, { 8'h1E}, { 8'h30}, { 8'h1F}, { 8'h00}}; // s
			8'h74: data <= {{8'h08}, { 8'h0C}, { 8'h3E}, { 8'h0C}, { 8'h0C}, { 8'h2C}, { 8'h18}, { 8'h00}}; // t
			8'h75: data <= {{8'h00}, { 8'h00}, { 8'h33}, { 8'h33}, { 8'h33}, { 8'h33}, { 8'h6E}, { 8'h00}}; // u
			8'h76: data <= {{8'h00}, { 8'h00}, { 8'h33}, { 8'h33}, { 8'h33}, { 8'h1E}, { 8'h0C}, { 8'h00}}; // v
			8'h77: data <= {{8'h00}, { 8'h00}, { 8'h63}, { 8'h6B}, { 8'h7F}, { 8'h7F}, { 8'h36}, { 8'h00}}; // w
			8'h78: data <= {{8'h00}, { 8'h00}, { 8'h63}, { 8'h36}, { 8'h1C}, { 8'h36}, { 8'h63}, { 8'h00}}; // x
			8'h79: data <= {{8'h00}, { 8'h00}, { 8'h33}, { 8'h33}, { 8'h33}, { 8'h3E}, { 8'h30}, { 8'h1F}}; // y
			8'h7A: data <= {{8'h00}, { 8'h00}, { 8'h3F}, { 8'h19}, { 8'h0C}, { 8'h26}, { 8'h3F}, { 8'h00}}; // z 
            
            default: data <= {{8'h00}, { 8'h00}, { 8'h00}, { 8'h00}, { 8'h00}, { 8'h00}, { 8'h00}, { 8'h00}}; // space
		endcase
	end

endmodule
